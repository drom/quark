module (/*AUTOARG*/);
/*AUTOINPUT*/
/*AUTOOUTPUT*/

/* let ir = input(); */
/* let irs = ir.splice(8); */
/* let pc = input(); */
/* let tailLength = ir.slice(8) */
/* let tailOffset =
*/

endmodule
