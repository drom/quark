
module imm (clk, reset_n, ti, te, to);
input           clk;
input           reset_n;
input           ti;
input           te;
output          to;

// declarations
always @(l0)
begin
l0
end

endmodule
